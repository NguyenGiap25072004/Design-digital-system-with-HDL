module NOT (
    input wire a_i,
    output wire y_o
);
assign y_o = ~a_i;

endmodule